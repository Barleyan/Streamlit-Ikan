��U      �sklearn.linear_model._base��LinearRegression���)��}�(�fit_intercept���copy_X���n_jobs�N�positive���n_features_in_�K�coef_��joblib.numpy_pickle��NumpyArrayWrapper���)��}�(�subclass��numpy��ndarray����shape�K���order��C��dtype�h�dtype����f8�����R�(K�<�NNNJ����J����K t�b�
allow_mmap���numpy_array_alignment_bytes�Kub���������������        �=�HcJA@�S�sa�X��h���A@�* �Zj%�c�RZ�E@��;��,%�9%6�A�:�-Α�>@�D}�����f��Q@��+��xE@�� �ӠE�T���nb@�\ǥ��O�F���@%YxQP�꿹!�Ķ%��!�^���g:����-@�_��/@�9       �rank_�K�	singular_�h)��}�(hhhK��hhhhh �h!Kub�����=҄(�@�M�N���@f� �k�@��M��o@Dj�/O\@j\��a�G@��nA@�|]��.@,�M�S)@p 앒@�-���7@8�3L?@�R$p��	@���K��?�M��[N�?��^���?��(�?���iMH�?_���rI�?jx{�0�?        �_       �
intercept_��numpy.core.multiarray��scalar���hC��F��Qf@���R��_sklearn_version��1.5.1�ub.